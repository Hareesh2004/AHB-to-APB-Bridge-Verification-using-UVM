package ahb2apb_pkg;

        import uvm_pkg::*;

        `include "uvm_macros.svh"

        `include "ahb_xtn.sv"
        `include "ahb_agent_config.sv"
        `include "apb_agent_config.sv"
        `include "ahb2apb_env_config.sv"

        `include "ahb_driver.sv"
        `include "ahb_monitor.sv"
        `include "ahb_sequencer.sv"
        `include "ahb_agent.sv"
        `include "ahb_agent_top.sv"
        `include "ahb_seqs.sv"

        `include "apb_xtn.sv"
        `include "apb_driver.sv"
        `include "apb_monitor.sv"
        `include "apb_sequencer.sv"
        `include "apb_agent.sv"
        `include "apb_agent_top.sv"

//      `include "ahb2apb_virtual_sequencer.sv"
//      `include "ahb2apb_virtual_seqs.sv"
        `include "ahb2apb_sb.sv"

        `include "ahb2apb_env.sv"
        `include "ahb2apb_test.sv"

endpackage

